`timescale 1ns / 1ps

module led_test (
                  clk,           // 开发板上输入时钟: 50Mhz
                  rst_n,         // 开发板上输入复位按键
                  led            // 输出LED灯,用于控制开发板上LED
             );
             
//===========================================================================
// PORT declarations
//===========================================================================
input clk;
input rst_n;
output led;

//寄存器定义
reg [31:0] timer;                  
reg led;


//===========================================================================
// 计数器计数:循环计数0~2秒
//===========================================================================
  always @(posedge clk or negedge rst_n)    //检测时钟的上升沿和复位的下降沿
    begin
      if (~rst_n)                           //复位信号低有效
          timer <= 0;                       //计数器清零
      else if (timer == 32'd99_999_999)     //开发板使用的晶振为50MHz，2秒计数(50M*2-1=99_999_999)
          timer <= 0;                       //计数器计到2秒，计数器清零
      else
		    timer <= timer + 1'b1;            //计数器加1
    end

//===========================================================================
// LED灯控制
//===========================================================================
  always @(posedge clk or negedge rst_n)   //检测时钟的上升沿和复位的下降沿
    begin
      if (~rst_n)                          //复位信号低有效
          led <= 1'b1;                  	 //LED灯输出为高
      else if (timer == 32'd49_999_999)    //计数器计到1秒，
          led <= 1'b0;                     //LED点亮
      else if (timer == 32'd99_999_999)    //计数器计到2秒，
          led <= 1'b1;                     //LED熄灭
    end
endmodule

