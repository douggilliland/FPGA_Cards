
module cv_altclkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
