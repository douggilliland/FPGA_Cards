
library ieee; 
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all; 
entity led_jt is 
port( 
      led_bit :out std_logic;                   --????????
      led_out :out std_logic_vector(7 downto 0) --????7???
    ); 
end led_jt ; 
architecture bhv of led_jt is 
begin  
  led_bit<= '0';             --?????????????
                             --????????

  led_out <="11111001";      --???????1??????
                             --?????7???????????????????
end bhv; 

