
module c10_altclkctrl (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
