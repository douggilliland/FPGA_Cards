// c10_altclkctrl.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module c10_altclkctrl (
		input  wire  inclk,  //  altclkctrl_input.inclk
		output wire  outclk  // altclkctrl_output.outclk
	);

	c10_altclkctrl_altclkctrl_0 altclkctrl_0 (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
